--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   16:53:58 10/28/2016
-- Design Name:   
-- Module Name:   D:/Arquitectura/Componentes/MUX4/tb_MUXF.vhd
-- Project Name:  MUX4
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: MUXF
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY tb_MUXF IS
END tb_MUXF;
 
ARCHITECTURE behavior OF tb_MUXF IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT MUXF
    PORT(
         A : IN  std_logic_vector(31 downto 0);
         B : IN  std_logic_vector(31 downto 0);
         C : IN  std_logic_vector(31 downto 0);
         D : IN  std_logic_vector(31 downto 0);
         Sc : IN  std_logic_vector(1 downto 0);
         S : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal A : std_logic_vector(31 downto 0) := (others => '0');
   signal B : std_logic_vector(31 downto 0) := (others => '0');
   signal C : std_logic_vector(31 downto 0) := (others => '0');
   signal D : std_logic_vector(31 downto 0) := (others => '0');
   signal Sc : std_logic_vector(1 downto 0) := (others => '0');

 	--Outputs
   signal S : std_logic_vector(31 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
  
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: MUXF PORT MAP (
          A => A,
          B => B,
          C => C,
          D => D,
          Sc => Sc,
          S => S
        ); 

   -- Stimulus process
   stim_proc: process
   begin		
		A <= "00000000000000000000000000000000";
		B <= "00000000000000000000000000000001";
		C <= "00000000000000000000000000000010";
		D <= "00000000000000000000000000000100";
		Sc <= "00";
		wait for 20 ns;
		Sc <= "01";
		wait for 20 ns;
		Sc <= "10";
		wait for 20 ns;
		Sc <= "11";
      wait;
   end process;

END;
